*
**********************************************************
*
* PDTC114EU
*
* NXP Semiconductors
*
* Resistor equipped NPN transistor (RET)
* IC   = 100 mA
* VCEO = 50 V
* hFE  = min. 30 @ 5V/5mA
* R1   = 10 Kohm
* R2   = 10 Kohm
*
*
* Package pinning does not match Spice model pinning.
* Package: SOT 323
*
* Package Pin 1: Base
* Package Pin 2: Emitter
* Package Pin 3: Collector
*
*
* Extraction date (week/year): 43/2014
* Simulator: Spice 3
*
**********************************************************
*sb#
* Please note: ---Resistances R1 and R2 are not part of the
* model and have to be added separately.---
* Diode D is dedicated to improve modeling in  reverse
* area of operation and does not reflect a physical device.
*
.SUBCKT PDTC114EU 1 2 3
*
Q1 1 4 3 MAIN
D1 2 1 DIODE
R1 2 4 10K
R2 4 3 10K
.MODEL MAIN NPN
+ IS = 7.342E-015
+ NF = 0.9765
+ ISE = 4.422E-015
+ NE = 1.742
+ BF = 296
+ IKF = 0.1257
+ VAF = 45.06
+ NR = 0.974
+ ISC = 8.521E-016
+ NC = 1.094
+ BR = 17.5
+ IKR = 1
+ VAR = 39
+ RB = 160
+ IRB = 0.000145
+ RBM = 4.2
+ RE = 0.3998
+ RC = 0.5587
+ XTB = 0
+ EG = 1.11
+ XTI = 3
+ CJE = 1.014E-011
+ VJE = 0.67
+ MJE = 0.3454
+ TF = 5.92E-010
+ XTF = 25
+ VTF = 2
+ ITF = 0.18
+ PTF = 0
+ CJC = 2.96E-012
+ VJC = 0.4591
+ MJC = 0.2956
+ XCJC = 1
+ TR = 8.7E-008
+ CJS = 0
+ VJS = 0.75
+ MJS = 0.333
+ FC = 0.78
.MODEL DIODE D
+ IS = 1.077E-015
+ N = 0.988
+ BV = 1000
+ IBV = 0.001
+ RS = 857.2
+ CJO = 0
+ VJ = 1
+ M = 0.5
+ FC = 0
+ TT = 0
+ EG = 1.11
+ XTI = 3
.ENDS
