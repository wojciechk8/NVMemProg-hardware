** Standard Linear Ics Macromodels, 1993.
** CONNECTIONS :
* 1 NON-INVERTING INPUT
* 2 INVERTING INPUT
* 3 POSITIVE POWER SUPPLY
* 4 NEGATIVE POWER SUPPLY
* 5 OUTPUT
.SUBCKT TS912 2 1 4 5 3
**********************************************************
.MODEL MDTH D IS=1E-8 KF=6.563355E-14 CJO=10F
* INPUT STAGE
CIP 2 5 1.500000E-12
CIN 1 5 1.500000E-12
EIP 10 5 2 5 1
EIN 16 5 1 5 1
RIP 10 11 6.500000E+00
RIN 15 16 6.500000E+00
RIS 11 15 7.655100E+00
DIP 11 12 MDTH 400E-12
DIN 15 14 MDTH 400E-12
VOFP 12 13 DC 0.000000E+00
VOFN 13 14 DC 0
IPOL 13 5 4.000000E-05
CPS 11 15 3.82E-08
DINN 17 13 MDTH 400E-12
VIN 17 5 -0.5000000e+00
DINR 15 18 MDTH 400E-12
VIP 4 18 -0.5000000E+00
FCP 4 5 VOFP 7.750000E+00
FCN 5 4 VOFN 7.750000E+00
* AMPLIFYING STAGE
FIP 5 19 VOFP 5.500000E+02
FIN 5 19 VOFN 5.500000E+02
RG1 19 5 5.087344E+05
RG2 19 4 5.087344E+05
CC 19 29 2.200000E-08
HZTP 30 29 VOFP 12.33E+02
HZTN  5 30 VOFN 12.33E+02
DOPM 19 22 MDTH 400E-12
DONM 21 19 MDTH 400E-12
HOPM 22 28 VOUT 3135
VIPM 28 4 150
HONM 21 27 VOUT 3135
VINM 5 27 150
EOUT 26 23 19 5 1
VOUT 23 5 0
ROUT 26 3 65
COUT 3 5 1.000000E-12
DOP 19 68 MDTH 400E-12
VOP 4 25 1.924
HSCP 68 25 VSCP1 1E8
DON 69 19 MDTH 400E-12
VON 24 5 2.4419107
HSCN 24 69 VSCN1 1.5E8
VSCTHP 60 61 0.1375
DSCP1 61 63 MDTH 400E-12
VSCP1 63 64 0
ISCP 64 0 1.000000E-8
DSCP2 0 64 MDTH 400E-12
DSCN2 0 74 MDTH 400E-12
ISCN 74 0 1.000000E-8
VSCN1 73 74 0
DSCN1 71 73 MDTH 400E-12
VSCTHN 71 70 -0.75
ESCP 60 0 2 1 500
ESCN 70 0 2 1 -2000
.ENDS
