*
**********************************************************
*
* BC807
*
* NXP Semiconductors
*
* General purpose PNP transistor
* IC   = 500 mA
* VCEO = 45 V 
* hFE  = 100 - 600 @ 1V/100mA
* 
*
*
*
* Package pinning does not match Spice model pinning.
* Package: SOT 23
* 
* Package Pin 1: Base
* Package Pin 2: Emitter
* Package Pin 3: Collector
* 
*
* 
* Simulator: Spice 2        
*
**********************************************************
*#
.MODEL QBC807 PNP 
+     IS=1.08E-13
+     NF=0.99
+     ISE=2.713E-14
+     NE=1.4
+     BF=385.7
+     IKF=0.3603
+     VAF=31.29
+     NR=0.9849
+     ISC=5.062E-13
+     NC=1.295
+     BR=20.57
+     IKR=0.054
+     VAR=11.62
+     RB=1
+     IRB=1E-06
+     RBM=0.5
+     RE=0.1415
+     RC=0.2623
+     XTB=0
+     EG=1.11
+     XTI=3
+     CJE=5.114E-11
+     VJE=0.8911
+     MJE=0.4417
+     TF=7.359E-10
+     XTF=1.859
+     VTF=3.813
+     ITF=0.4393
+     PTF=0
+     CJC=2.656E-11
+     VJC=0.62
+     MJC=0.4836
+     XCJC=0.459
+     TR=5.00E-08
+     CJS=0
+     VJS=0.75
+     MJS=0.333
+     FC=0.99
*##
*
